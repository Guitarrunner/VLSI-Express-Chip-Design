module sebas
